NOR_X1 Layout and Schematic Circuits

* Technology Dependent design rules/parameters
.include /CMC/setups/ensc450/HSPICE/cmosp18/rules.inc
* Wm#, Awd# parameters etc. all specified in the rules.inc file above

* Transistor models 
.protect
.LIB `/CMC/setups/ensc450/HSPICE/cmosp18/log018.l' SS  $ typical process corner.
.unprotect
* WORST CASE SIMULATION

* Supply Sources
.param pwr=1.05 
.temp 125
Vvdd  VDD!  0 dc pwr
Vgnd  GND!  0 dc 0

* Schematic Logic
MNMOS3 Z_S B GND! GND!  NCH  L=180E-9 W=500E-9 AD=+2.40000000E-13 AS=+2.40000000E-13
+PD=+1.09600000E-05 PS=+1.09600000E-05 NRD=+5.40000000E-01 NRS=+5.40000000E-01
+M=1.0
MNMOS2 Z_S A GND! GND!  NCH  L=180E-9 W=500E-9 AD=+2.40000000E-13 AS=+2.40000000E-13
+PD=+1.09600000E-05 PS=+1.09600000E-05 NRD=+5.40000000E-01 NRS=+5.40000000E-01
+M=1.0
MPMOS1 Z_S B NET036 VDD!  PCH  L=180E-9 W=2E-6 AD=+9.60000000E-13 AS=+9.60000000E-13
+PD=+4.96000000E-06 PS=+4.96000000E-06 NRD=+1.35000000E-01 NRS=+1.35000000E-01
+M=1.0
MPMOS0 NET036 A VDD! VDD!  PCH  L=180E-9 W=2E-6 AD=+9.60000000E-13
+AS=+9.60000000E-13 PD=+4.96000000E-06 PS=+4.96000000E-06 NRD=+1.35000000E-01
+NRS=+1.35000000E-01 M=1.0

* Extracted Layout Logic
MPMOS3 VDD! A 1 VDD!  PCH  L=180.000000682412E-9 W=1.99999999495049E-6
+AD=959.999983153603E-15 AS=540.000010852693E-15 PD=2.96000007438124E-6
+PS=539.999973625527E-9 NRD=+1.35000034E-01 NRS=+1.35000000E-01 M=1.0
MPMOS4 1 B Z_E VDD!  PCH  L=180.000000682412E-9 W=1.99999999495049E-6
+AD=540.000010852693E-15 AS=959.999983153603E-15 PD=539.999973625527E-9
+PS=2.96000007438124E-6 NRD=+1.35000000E-01 NRS=+1.35000034E-01 M=1.0
MNMOS5 GND! A Z_E GND!  NCH  L=180.000000682412E-9 W=499.999998737621E-9
+AD=239.999995788401E-15 AS=135.000002713173E-15 PD=1.46000002132496E-6
+PS=539.999973625527E-9 NRD=+5.40000028E-01 NRS=+5.40000001E-01 M=1.0
MNMOS6 Z_E B GND! GND!  NCH  L=180.000000682412E-9 W=499.999998737621E-9
+AD=135.000002713173E-15 AS=239.999995788401E-15 PD=539.999973625527E-9
+PS=1.46000002132496E-6 NRD=+5.40000001E-01 NRS=+5.40000028E-01 M=1.0 

Cload_S Z_S 0 load
Cload_E Z_E 0 load

* Input Stimuli (Step response)
VB  B  0 PWL(0n 0 5ns 0 6ns 0 11ns 0 12ns 0 17ns 0 19ns 0 23ns 0)
VA  A  0 PWL(0n pwr 3ns pwr 4ns 0 8ns 0  9ns pwr 13ns pwr 15ns 0 19ns 0 21ns pwr 23ns pwr)

* Simulation Parameters ************************ 
.tran 0.01ps 25ns START=0 sweep load POI 2 2fF 10fF 

.graph V(A)
.graph V(B)
.graph V(Z_S)
.graph V(Z_E)
.option post
************************************************
* Various Timing Measurements 

* Measure propogation delay from rising edge of input A to falling edge of output Z
.meas tran tpdf_1ns      trig v(A) val='pwr*0.5' cross=2
+                        targ v(Z_E) val='pwr*0.5' cross=2 
.meas tran tpdf_2ns      trig v(A) val='pwr*0.5' cross=4
+                        targ v(Z_E) val='pwr*0.5' cross=4

* Rise propogation delay
.meas tran tpdr_1ns      trig v(A) val='pwr*0.5' cross=1
+                        targ v(Z_E) val='pwr*0.5' cross=1 
.meas tran tpdr_2ns      trig v(A) val='pwr*0.5' cross=3
+			 targ v(Z_E) val='pwr*0.5' cross=3

* Rise Time
.meas tran ttr_1ns       trig v(Z_E) val='pwr*0.2' rise=1
+                        targ v(Z_E) val='pwr*0.8' rise=1
.meas tran ttr_2ns       trig v(Z_E) val='pwr*0.2' rise=2
+                        targ v(Z_E) val='pwr*0.8' rise=2

* Fall Time
.meas tran ttf_1ns       trig v(Z_E) val='pwr*0.8' fall=1
+                        targ v(Z_E) val='pwr*0.2' fall=1
.meas tran ttf_2ns       trig v(Z_E) val='pwr*0.8' fall=2
+                        targ v(Z_E) val='pwr*0.2' fall=2

************************************************
.end
  
