NOR_X1 Layout Schematic

* Technology Dependent design rules/parameters
.include /CMC/setups/ensc450/HSPICE/cmosp18/rules.inc
* Wm#, Awd# parameters etc. all specified in the rules.inc file above

* Transistor models 
.protect
.LIB `/CMC/setups/ensc450/HSPICE/cmosp18/log018.l' SS  $ typical process corner.
.unprotect
* WORST CASE SIMULATION

* Supply Sources
.param pwr=1.05 
.temp 125
Vvdd  VDD!  0 dc pwr
Vgnd  GND!  0 dc 0

* Logic 
MNMOS3 VDD! B 1 VDD!  PCH  L=180.000000682412E-9 W=3.99999998990097E-6
+AD=1.91999996630721E-12 AS=1.08000002170539E-12 PD=4.95999984195805E-6
+PS=539.999973625527E-9 NRD=+6.75000002E-02 NRS=+6.75000002E-02 M=1.0
MNMOS4 1 A Z VDD!  PCH  L=180.000000682412E-9 W=3.99999998990097E-6
+AD=1.08000002170539E-12 AS=1.91999996630721E-12 PD=539.999973625527E-9
+PS=4.95999984195805E-6 NRD=+6.75000002E-02 NRS=+6.75000002E-02 M=1.0
MPMOS5 GND! B Z GND!  NCH  L=180.000000682412E-9 W=999.999997475243E-9
+AD=479.999991576802E-15 AS=270.000005426346E-15 PD=1.95999996321916E-6
+PS=539.999973625527E-9 NRD=+2.70000014E-01 NRS=+2.70000001E-01 M=1.0
MPMOS6 Z A GND! GND!  NCH  L=180.000000682412E-9 W=999.999997475243E-9
+AD=270.000005426346E-15 AS=479.999991576802E-15 PD=539.999973625527E-9
+PS=1.95999996321916E-6 NRD=+2.70000001E-01 NRS=+2.70000014E-01 M=1.0

Cload z 0 load

* Input Stimuli (Step response)
VB  b  0 PWL(0n 0 5ns 0 6ns 0 11ns 0 12ns 0 17ns 0 19ns 0 23ns 0)
VA  a  0 PWL(0n pwr 3ns pwr 4ns 0 8ns 0  9ns pwr 13ns pwr 15ns 0 19ns 0 21ns pwr 23ns pwr)

* Simulation Parameters ************************ 
.tran 0.01ps 25ns START=0 sweep load POI 2 2fF 10fF 

.graph V(a)
.graph V(b)
.graph V(z)
.option post
************************************************
* Various Timing Measurements 

* Measure propogation delay from rising edge of input A to falling edge of output Z
.meas tran tpdf_1ns      trig v(a) val='pwr*0.5' cross=2
+                        targ v(z) val='pwr*0.5' cross=2 
.meas tran tpdf_2ns      trig v(a) val='pwr*0.5' cross=4
+                        targ v(z) val='pwr*0.5' cross=4

* Rise propogation delay
.meas tran tpdr_1ns      trig v(a) val='pwr*0.5' cross=1
+                        targ v(z) val='pwr*0.5' cross=1 
.meas tran tpdr_2ns      trig v(a) val='pwr*0.5' cross=3
+			 targ v(z) val='pwr*0.5' cross=3

* Rise Time
.meas tran ttr_1ns       trig v(z) val='pwr*0.2' rise=1
+                        targ v(z) val='pwr*0.8' rise=1
.meas tran ttr_2ns       trig v(z) val='pwr*0.2' rise=2
+                        targ v(z) val='pwr*0.8' rise=2

* Fall Time
.meas tran ttf_1ns       trig v(z) val='pwr*0.8' fall=1
+                        targ v(z) val='pwr*0.2' fall=1
.meas tran ttf_2ns       trig v(z) val='pwr*0.8' fall=2
+                        targ v(z) val='pwr*0.2' fall=2

************************************************
.end
  
