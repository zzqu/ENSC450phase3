NOR_X1_L3

* Technology Dependent design rules/parameters
.include /CMC/setups/ensc450/HSPICE/cmosp18/rules.inc
* Wm#, Awd# parameters etc. all specified in the rules.inc file above

* Transistor models 
.protect
.LIB `/CMC/setups/ensc450/HSPICE/cmosp18/log018.l' SS  $ typical process corner.
.unprotect
* WORST CASE SIMULATION

* Supply Sources
.param pwr=1.05 
.temp 125
Vvdd  VDD!  0 dc pwr
Vgnd  GND!  0 dc 0

* Logic 
MNMOS3 Z B GND! GND!  NCH  L=180E-9 W=1E-6 AD=+4.80000000E-13 AS=+4.80000000E-13
+PD=+2.96000000E-06 PS=+2.96000000E-06 NRD=+2.70000000E-01 NRS=+2.70000000E-01
+M=1.0
MNMOS2 Z A GND! GND!  NCH  L=180E-9 W=1E-6 AD=+4.80000000E-13 AS=+4.80000000E-13
+PD=+2.96000000E-06 PS=+2.96000000E-06 NRD=+2.70000000E-01 NRS=+2.70000000E-01
+M=1.0
MPMOS1 Z B NET15 NET15  PCH  L=180E-9 W=4E-6 AD=+1.92000000E-12 AS=+1.92000000E-12
+PD=+8.96000000E-06 PS=+8.96000000E-06 NRD=+6.75000000E-02 NRS=+6.75000000E-02
+M=1.0
MPMOS0 NET15 A VDD! VDD!  PCH  L=180E-9 W=4E-6 AD=+1.92000000E-12
+AS=+1.92000000E-12 PD=+8.96000000E-06 PS=+8.96000000E-06 NRD=+6.75000000E-02
+NRS=+6.75000000E-02 M=1.0

Cload z 0 load

* Input Stimuli (Step response)
VB  b  0 PWL(0n 0 5ns 0 6ns 0 11ns 0 12ns 0 17ns 0 19ns 0 23ns 0)
VA  a  0 PWL(0n pwr 3ns pwr 4ns 0 8ns 0  9ns pwr 13ns pwr 15ns 0 19ns 0 21ns pwr 23ns pwr)

* Simulation Parameters ************************ 
.tran 0.01ps 25ns START=0 sweep load POI 2 2fF 10fF 

.graph V(a)
.graph V(b)
.graph V(z)
.option post
************************************************

.end
  
